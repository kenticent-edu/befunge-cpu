----------------------------------------------------------------------------------
-- Company:
-- Engineer:
--
-- Create Date: 03/16/2021 06:09:57 PM
-- Design Name:
-- Module Name: rom_64x16 - Behavioral
-- Project Name:
-- Target Devices:
-- Tool Versions:
-- Description:
--
-- Dependencies:
--
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
----------------------------------------------------------------------------------


library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity rom_64x16 is
port (
address  : in STD_LOGIC_VECTOR (5 downto 0);
clk      : in STD_LOGIC;
data_out : out STD_LOGIC_VECTOR (15 downto 0)
);
end entity;

architecture rom_64x16_arch of rom_64x16 is

type ROM_type is array ( 0 to 63 ) of std_logic_vector(15 downto 0);

constant ROM : ROM_type := ( 0 => "0000010001110101",
1 => "0010100100001101",
2 => "0011110000110110",
3 => "0101000111001100",
4 => "1111001000000011",
5 => "1111101100000011",
6 => "0001000110101100",
7 => "0010101100001010",
8 => "1001111111111101",
9 => "1000110010110010",
10 => "1010100111001001",
11 => "0100110100111110",
12 => "0101010001110010",
13 => "0001011100111010",
14 => "1011111100100011",
15 => "0001111011110011",
16 => "1001000010001010",
17 => "0001010011101111",
18 => "1010100000101001",
19 => "1011111000000111",
20 => "1111111001100100",
21 => "0111111011101111",
22 => "0111011110011101",
23 => "1011100001011011",
24 => "1111010011010000",
25 => "1001111010000110",
26 => "1111100001110011",
27 => "1010011010010011",
28 => "0001110001001100",
29 => "0100111111010000",
30 => "0111101010001000",
31 => "1111100111110010",
32 => "1001001010001111",
33 => "0100101010001111",
34 => "0010101100000110",
35 => "1101000001001110",
36 => "0100010100010100",
37 => "1101011011100101",
38 => "1111011001111010",
39 => "0010110111101000",
40 => "1110001001101100",
41 => "1110010111000101",
42 => "1100110110001110",
43 => "0010111110100111",
44 => "1001110111011011",
45 => "1010100100001000",
46 => "0011100001111100",
47 => "1011110010011000",
48 => "0011000011011000",
49 => "1000110100111100",
50 => "1100001100001111",
51 => "0101110111011001",
52 => "1110100100100111",
53 => "0011100010011011",
54 => "1010101000001001",
55 => "0101001110000011",
56 => "0011001011011010",
57 => "0101000100101100",
58 => "0000110000001100",
59 => "1111011101001001",
60 => "0001011111010000",
61 => "0111010110100110",
62 => "1101011000111110",
63 => "0111110111000001");

begin

process(clk)
begin
            if clk'event and clk = '1' then
                data_out <= ROM (to_integer(unsigned(address)));
            end if;
end process;
end architecture;